






// post process / activation 

// simple post process

// integer 