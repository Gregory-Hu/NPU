














// ----------------------------------------------------------
// SOC Interface 
//     - APB Command interface 
//     - AXI (dedicated memory bandwidth)
//     - local mmu
//     - CHI Stash
//     - interrupt


// ----------------------------------------------------------
// Scratch SRAM


// ----------------------------------------------------------
// NPU AI Engine (Matrix computation)
//     - MAC Array
//     - activation unit 
//     - Load Store Unit
//     - Transpose Unit (Pre Post)


// ----------------------------------------------------------
// USC_RVV Cores
//     - Post Process Vector Computation
//     - branching flow control
//     - streaming vector processor 


// ----------------------------------------------------------
// Shared Cache
//     - time locality data


// ----------------------------------------------------------
// do we need hts to dynamicly schedule work load 

