

module npu_fast_post_process #(
) ( 
  input wire clk, 
  input wire reset_n,

  // NN Data Stream

  // Processed Result
)

endmodule 